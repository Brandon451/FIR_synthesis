//Transpose form

module fir4rca #(
    parameter w = 16
)(
    input clk,
    input reset,
    input [w-1:0] a,
    output logic [w+1:0] s
);

//Pipeline for inputs
logic [w-1:0] ar;

//Pipeline for sums
logic [w:0]     sum1;
logic [w:0]     sum1r;
logic [w+1:0]   sum2;
logic [w+1:0]   sum2r;
logic [w+1:0]   sum3;

logic [w-1:0]   rca1_s;
logic [w:0]     rca2_s;
logic [w+1:0]   rca3_s;
logic [w:0]     cr2;
logic [w+1:0]   dr3;
logic [w:0]     rca1_co;    //Carry in
logic [w+1:0]   rca2_co;
logic [w+2:0]   rca3_co;

logic [w+1:0]   sum;

always_comb begin
    rca1_co[0] = 0;
    for (int i=0; i<w; i++)
        {rca1_co[i+1], rca1_s[i]} = ar[i] + a[i] + rca1_co[i];
    sum1 = {rca1_co[w], rca1_s};
end

always_comb begin
    rca2_co[0] = 0;
    cr2 = {1'b0,a};
    for(int i=0; i<w+1; i++)
        {rca2_co[i+1],rca2_s[i]} = sum1r[i] + cr2[i] + rca2_co[i];
    sum2 = {rca2_co[w+1],rca2_s};
end

always_comb begin    
    rca3_co[0] = 0;
    dr3 = {2'b0,a};
    for(int i=0; i<w+2; i++)
        {rca3_co[i+1],rca3_s[i]} = sum2r[i] + dr3[i] + rca3_co[i];
end

always_comb
    sum = rca3_s;

//Shift register to store outputs
always_ff @(posedge clk)			// or just always -- always_ff tells tools you intend D flip flops
    if(reset) begin					// reset forces all registers to 0 for clean start of test
        ar <= 'b0;
        sum1r <= 'b0;
        sum2r <= 'b0;
        s  <= 'b0;
    end
    else begin					    // normal operation -- Dffs update on posedge clk
        ar <= a;
        sum1r <= sum1;
        sum2r <= sum2;
        s  <= sum; 
    end

endmodule